`define wTime10 5'd00
`define wTime11 5'd03
`define wTime12 5'd06
`define wTime13 5'd09
`define wTime14 5'd12
`define wTime15 5'd15
`define wTime16 5'd18
`define wTime17 5'd21
`define wTime20 5'd00
`define wTime21 5'd03
`define wTime22 5'd04
`define wTime23 5'd06
`define wTime24 5'd04
`define wTime25 5'd09
`define wTime26 5'd10
`define wTime27 5'd12
`define wTime30 5'd00
`define wTime31 5'd03
`define wTime32 5'd04
`define wTime33 5'd05
`define wTime34 5'd06
`define wTime35 5'd07
`define wTime36 5'd08
`define wTime37 5'd09